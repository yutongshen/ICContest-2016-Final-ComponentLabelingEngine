
module CLE_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
  CLKINVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module CLE_DW01_inc_1 ( A, SUM );
  input [10:0] A;
  output [10:0] SUM;

  wire   [10:2] carry;

  ADDHXL U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADDHXL U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(carry[10]), .B(A[10]), .Y(SUM[10]) );
  CLKINVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module CLE_DW01_inc_2 ( A, SUM );
  input [10:0] A;
  output [10:0] SUM;
  wire   n1;
  wire   [10:2] carry;

  ADDHXL U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHXL U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  CLKINVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  CLKINVX1 U2 ( .A(SUM[0]), .Y(n1) );
  XOR2X1 U3 ( .A(carry[10]), .B(A[10]), .Y(SUM[10]) );
endmodule


module CLE_DW01_inc_3 ( A, SUM );
  input [20:0] A;
  output [20:0] SUM;

  wire   [20:2] carry;

  ADDHXL U1_1_19 ( .A(A[19]), .B(carry[19]), .CO(carry[20]), .S(SUM[19]) );
  ADDHXL U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  ADDHXL U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  ADDHXL U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  ADDHXL U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  ADDHXL U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  ADDHXL U1_1_15 ( .A(A[15]), .B(carry[15]), .CO(carry[16]), .S(SUM[15]) );
  ADDHXL U1_1_17 ( .A(A[17]), .B(carry[17]), .CO(carry[18]), .S(SUM[17]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_16 ( .A(A[16]), .B(carry[16]), .CO(carry[17]), .S(SUM[16]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_18 ( .A(A[18]), .B(carry[18]), .CO(carry[19]), .S(SUM[18]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHXL U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADDHXL U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  XOR2XL U1 ( .A(carry[20]), .B(A[20]), .Y(SUM[20]) );
  INVXL U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module CLE ( clk, reset, rom_q, rom_a, sram_q, sram_a, sram_d, sram_wen, 
        finish );
  input [7:0] rom_q;
  output [6:0] rom_a;
  input [7:0] sram_q;
  output [9:0] sram_a;
  output [7:0] sram_d;
  input clk, reset;
  output sram_wen, finish;
  wire   n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, index_buffer_28__7_, index_buffer_28__6_, index_buffer_28__5_,
         index_buffer_28__4_, index_buffer_28__3_, index_buffer_28__2_,
         index_buffer_28__1_, index_buffer_28__0_, index_buffer_29__6_,
         index_buffer_29__4_, index_buffer_29__2_, index_buffer_29__0_, rw,
         rd_sram, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79,
         N80, N81, N82, N83, N84, N85, N86, N87, N88, N114, N115, N116, N117,
         N118, N119, N120, N121, N122, N123, N124, N138, N139, N140, N141,
         N142, N143, N144, N145, N146, N147, N148, N149, N150, N151, N152,
         N153, N154, N155, N156, N157, N158, N160, N161, N162, N163, N164,
         N165, N166, N168, N181, N182, N183, cs, N336, N337, N338, N339, N340,
         N341, N342, N343, N397, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n680,
         n690, n700, n710, n720, n730, n740, n7500, n7600, n7700, n7800, n7900,
         n8000, n8100, n820, n830, n840, n850, n860, n870, n880, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n11400, n1150,
         n1160, n1170, n11800, n11900, n12000, n12100, n12200, n12300, n12400,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n13800, n13900, n14000, n14100, n14210, n14340, n1440,
         n1450, n1460, n1470, n1480, n1490, n1500, n1510, n1520, n1530, n1540,
         n1550, n1560, n1570, n1580, n159, n1600, n1610, n1620, n1630, n1640,
         n1650, n1660, n167, n1680, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n1810, n1820, n1830, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n314,
         n326, n365, n366, n367, n368, n369, n370, n371, n372, n597, n599,
         n600, n601, n602, n603, n604, n606, n608, n610, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n707, n747, n748, n749, n7501, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n7601, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n7701, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n7801, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n7901, n791, n792, n793, n794, n795, n796, n797, n798, n799, n8001,
         n801, n802, n807, n808, n809, n8101, n811, n812, n813, n815, n818,
         n821, n1567, n826, n828, n923, n925, n927, n929, n931, n933, n935,
         n937, n941, n942, n943, n944, n945, n946, n947, n1134, n1135, n1136,
         n1137, n1138, n1139, n11401, n1141, n1142, n1143, n1144, n1175, n1176,
         n1177, n1178, n1179, n11801, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n11901, n1192, n1194, n1196, n1198, n1199,
         n12001, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n12101, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n12201, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n12301, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n12401, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n13801, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n13901, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n14001, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n14101, n1411, n1412, n14341, n1436, n1437, n1438;
  wire   [3:0] cnt;
  wire   [40:1] rd_buffer;
  wire   [7:0] index_cnt;
  wire   [20:0] times;
  wire   [4:0] rom_a_high;
  wire   [1:0] rom_a_low;
  wire   [4:0] read_addr_high;
  wire   [4:0] read_addr_low;
  wire   [4:0] write_addr_high;
  wire   [4:1] write_addr_low;
  wire   [2:0] re_cs;
  wire   [9:3] add_95_carry;

  EDFFTRX1 index_cnt_reg_7_ ( .RN(n1196), .D(N343), .E(n1412), .CK(clk), .Q(
        index_cnt[7]), .QN(n365) );
  EDFFTRX1 rd_buffer_reg_38_ ( .RN(n1196), .D(n238), .E(n1221), .CK(clk), .Q(
        n1241), .QN(n326) );
  EDFFTRX1 rd_buffer_reg_39_ ( .RN(n1196), .D(n1241), .E(n1221), .CK(clk), .Q(
        rd_buffer[39]), .QN(n1409) );
  EDFFTRX1 rd_buffer_reg_8_ ( .RN(n1198), .D(rd_buffer[7]), .E(n1221), .CK(clk), .Q(rd_buffer[8]), .QN(n1408) );
  EDFFTRX1 index_cnt_reg_1_ ( .RN(n1196), .D(N337), .E(n1412), .CK(clk), .Q(
        index_cnt[1]), .QN(n371) );
  EDFFTRX1 index_cnt_reg_2_ ( .RN(n1196), .D(N338), .E(n1412), .CK(clk), .Q(
        index_cnt[2]), .QN(n370) );
  EDFFTRX1 index_cnt_reg_3_ ( .RN(n1196), .D(N339), .E(n1412), .CK(clk), .Q(
        index_cnt[3]), .QN(n369) );
  EDFFTRX1 index_cnt_reg_4_ ( .RN(n1196), .D(N340), .E(n1412), .CK(clk), .Q(
        index_cnt[4]), .QN(n368) );
  EDFFTRX1 index_cnt_reg_5_ ( .RN(n1196), .D(N341), .E(n1412), .CK(clk), .Q(
        index_cnt[5]), .QN(n367) );
  EDFFTRX1 index_cnt_reg_6_ ( .RN(n1196), .D(N342), .E(n1412), .CK(clk), .Q(
        index_cnt[6]), .QN(n366) );
  EDFFTRX1 index_cnt_reg_0_ ( .RN(n1196), .D(N336), .E(n1412), .CK(clk), .Q(
        index_cnt[0]), .QN(n372) );
  EDFFTRX1 rd_sram_reg ( .RN(n1199), .D(1'b1), .E(n707), .CK(clk), .Q(rd_sram)
         );
  DFFTRX1 cnt_reg_3_ ( .D(N117), .RN(n1187), .CK(clk), .Q(cnt[3]) );
  DFFTRX1 cnt_reg_1_ ( .D(N115), .RN(n1187), .CK(clk), .Q(cnt[1]) );
  DFFTRX1 cnt_reg_2_ ( .D(N116), .RN(n1187), .CK(clk), .Q(cnt[2]) );
  DFFTRX1 read_addr_low_reg_1_ ( .D(N150), .RN(n1188), .CK(clk), .Q(
        read_addr_low[1]) );
  DFFTRX1 read_addr_low_reg_2_ ( .D(N151), .RN(n1188), .CK(clk), .Q(
        read_addr_low[2]) );
  DFFTRX1 read_addr_high_reg_1_ ( .D(N155), .RN(n1188), .CK(clk), .Q(
        read_addr_high[1]) );
  DFFTRX1 read_addr_low_reg_0_ ( .D(N149), .RN(n1188), .CK(clk), .Q(
        read_addr_low[0]) );
  DFFTRX1 read_addr_high_reg_0_ ( .D(N154), .RN(n1188), .CK(clk), .Q(
        read_addr_high[0]) );
  DFFTRX1 read_addr_high_reg_2_ ( .D(N156), .RN(n1188), .CK(clk), .Q(
        read_addr_high[2]) );
  DFFTRX1 read_addr_high_reg_3_ ( .D(N157), .RN(n1188), .CK(clk), .Q(
        read_addr_high[3]) );
  DFFTRX1 read_addr_high_reg_4_ ( .D(N158), .RN(n1188), .CK(clk), .Q(
        read_addr_high[4]) );
  DFFTRX1 write_addr_high_reg_0_ ( .D(N144), .RN(n1188), .CK(clk), .Q(
        write_addr_high[0]), .QN(n1242) );
  EDFFTRX1 times_reg_11_ ( .RN(n1199), .D(N79), .E(n1184), .CK(clk), .Q(
        times[11]), .QN(n1247) );
  EDFFTRX1 times_reg_14_ ( .RN(n1199), .D(N82), .E(n1184), .CK(clk), .Q(
        times[14]), .QN(n1244) );
  EDFFTRX1 times_reg_10_ ( .RN(n1199), .D(N78), .E(n1184), .CK(clk), .Q(
        times[10]), .QN(n1248) );
  EDFFTRX1 times_reg_13_ ( .RN(n1199), .D(N81), .E(n1184), .CK(clk), .Q(
        times[13]), .QN(n1245) );
  EDFFTRX1 times_reg_12_ ( .RN(n1199), .D(N80), .E(n1184), .CK(clk), .Q(
        times[12]), .QN(n1246) );
  EDFFTRX1 times_reg_20_ ( .RN(n1199), .D(N88), .E(n1184), .CK(clk), .Q(
        times[20]) );
  DFFTRX1 rom_a_high_reg_4_ ( .D(N124), .RN(n1187), .CK(clk), .Q(rom_a_high[4]) );
  EDFFTRX1 times_reg_15_ ( .RN(n1199), .D(N83), .E(n1184), .CK(clk), .Q(
        times[15]) );
  EDFFTRX1 times_reg_17_ ( .RN(n1199), .D(N85), .E(n1184), .CK(clk), .Q(
        times[17]) );
  EDFFTRX1 times_reg_1_ ( .RN(n12001), .D(N69), .E(n1184), .CK(clk), .Q(
        times[1]) );
  EDFFTRX1 times_reg_2_ ( .RN(n12001), .D(N70), .E(n1184), .CK(clk), .Q(
        times[2]) );
  EDFFTRX1 times_reg_16_ ( .RN(n1199), .D(N84), .E(n1184), .CK(clk), .Q(
        times[16]) );
  EDFFTRX1 times_reg_18_ ( .RN(n1199), .D(N86), .E(n1184), .CK(clk), .Q(
        times[18]) );
  EDFFTRX1 times_reg_4_ ( .RN(n12001), .D(N72), .E(n1184), .CK(clk), .Q(
        times[4]) );
  EDFFTRX1 times_reg_7_ ( .RN(n12001), .D(N75), .E(n1184), .CK(clk), .Q(
        times[7]) );
  EDFFTRX1 times_reg_19_ ( .RN(n1199), .D(N87), .E(n1184), .CK(clk), .Q(
        times[19]) );
  EDFFTRX1 times_reg_5_ ( .RN(n12001), .D(N73), .E(n1184), .CK(clk), .Q(
        times[5]) );
  EDFFTRX1 times_reg_8_ ( .RN(n1199), .D(N76), .E(n1184), .CK(clk), .Q(
        times[8]) );
  EDFFTRX1 times_reg_3_ ( .RN(n12001), .D(N71), .E(n1184), .CK(clk), .Q(
        times[3]) );
  EDFFTRX1 times_reg_6_ ( .RN(n12001), .D(N74), .E(n1184), .CK(clk), .Q(
        times[6]) );
  EDFFTRX1 times_reg_9_ ( .RN(n1199), .D(N77), .E(n1184), .CK(clk), .Q(
        times[9]) );
  EDFFTRX1 times_reg_0_ ( .RN(n12001), .D(N68), .E(n1184), .CK(clk), .Q(
        times[0]) );
  DFFTRX1 rom_a_high_reg_0_ ( .D(N120), .RN(n1187), .CK(clk), .Q(rom_a_high[0]) );
  DFFTRX1 rom_a_low_reg_1_ ( .D(N119), .RN(n1187), .CK(clk), .Q(rom_a_low[1])
         );
  DFFTRX1 rom_a_high_reg_1_ ( .D(N121), .RN(n1187), .CK(clk), .Q(rom_a_high[1]) );
  DFFTRX1 rom_a_high_reg_2_ ( .D(N122), .RN(n1187), .CK(clk), .Q(rom_a_high[2]) );
  DFFTRX1 rom_a_high_reg_3_ ( .D(N123), .RN(n1187), .CK(clk), .Q(rom_a_high[3]) );
  EDFFTRX1 index_buffer_reg_6__6_ ( .RN(n1206), .D(n106), .E(n11801), .CK(clk), 
        .Q(n105) );
  EDFFTRX1 index_buffer_reg_5__6_ ( .RN(n1206), .D(n105), .E(n1178), .CK(clk), 
        .Q(n104) );
  EDFFTRX1 index_buffer_reg_4__6_ ( .RN(n1206), .D(n104), .E(n1179), .CK(clk), 
        .Q(n103) );
  EDFFTRX1 index_buffer_reg_3__6_ ( .RN(n1206), .D(n103), .E(n11801), .CK(clk), 
        .Q(n102) );
  EDFFTRX1 index_buffer_reg_2__6_ ( .RN(n1206), .D(n102), .E(n1178), .CK(clk), 
        .Q(n101) );
  EDFFTRX1 index_buffer_reg_1__6_ ( .RN(n1206), .D(n101), .E(n1179), .CK(clk), 
        .Q(n100) );
  EDFFTRX1 index_buffer_reg_18__5_ ( .RN(n1205), .D(n91), .E(n1178), .CK(clk), 
        .Q(n90) );
  EDFFTRX1 index_buffer_reg_17__5_ ( .RN(n1205), .D(n90), .E(n1179), .CK(clk), 
        .Q(n89) );
  EDFFTRX1 index_buffer_reg_16__5_ ( .RN(n1205), .D(n89), .E(n11801), .CK(clk), 
        .Q(n880) );
  EDFFTRX1 index_buffer_reg_15__5_ ( .RN(n1205), .D(n880), .E(n1178), .CK(clk), 
        .Q(n870) );
  EDFFTRX1 index_buffer_reg_14__5_ ( .RN(n1205), .D(n870), .E(n1179), .CK(clk), 
        .Q(n860) );
  EDFFTRX1 index_buffer_reg_13__5_ ( .RN(n1205), .D(n860), .E(n11801), .CK(clk), .Q(n850) );
  EDFFTRX1 index_buffer_reg_12__5_ ( .RN(n1205), .D(n850), .E(n1178), .CK(clk), 
        .Q(n840) );
  EDFFTRX1 index_buffer_reg_11__5_ ( .RN(n1205), .D(n840), .E(n1179), .CK(clk), 
        .Q(n830) );
  EDFFTRX1 index_buffer_reg_10__5_ ( .RN(n1205), .D(n830), .E(n11801), .CK(clk), .Q(n820) );
  EDFFTRX1 index_buffer_reg_9__5_ ( .RN(n1205), .D(n820), .E(n1219), .CK(clk), 
        .Q(n8100) );
  EDFFTRX1 index_buffer_reg_8__5_ ( .RN(n1205), .D(n8100), .E(n12201), .CK(clk), .Q(n8000) );
  EDFFTRX1 index_buffer_reg_7__5_ ( .RN(n1204), .D(n8000), .E(n12201), .CK(clk), .Q(n7900) );
  EDFFTRX1 index_buffer_reg_6__5_ ( .RN(n1204), .D(n7900), .E(n1219), .CK(clk), 
        .Q(n7800) );
  EDFFTRX1 index_buffer_reg_5__5_ ( .RN(n1204), .D(n7800), .E(n1219), .CK(clk), 
        .Q(n7700) );
  EDFFTRX1 index_buffer_reg_4__5_ ( .RN(n1204), .D(n7700), .E(n12201), .CK(clk), .Q(n7600) );
  EDFFTRX1 index_buffer_reg_3__5_ ( .RN(n1204), .D(n7600), .E(n12201), .CK(clk), .Q(n7500) );
  EDFFTRX1 index_buffer_reg_2__5_ ( .RN(n1204), .D(n7500), .E(n1219), .CK(clk), 
        .Q(n740) );
  EDFFTRX1 index_buffer_reg_1__5_ ( .RN(n1204), .D(n740), .E(n1219), .CK(clk), 
        .Q(n730) );
  EDFFTRX1 index_buffer_reg_18__4_ ( .RN(n1203), .D(n64), .E(n12201), .CK(clk), 
        .Q(n63) );
  EDFFTRX1 index_buffer_reg_17__4_ ( .RN(n1203), .D(n63), .E(n1219), .CK(clk), 
        .Q(n62) );
  EDFFTRX1 index_buffer_reg_16__4_ ( .RN(n1203), .D(n62), .E(n1177), .CK(clk), 
        .Q(n61) );
  EDFFTRX1 index_buffer_reg_15__4_ ( .RN(n1203), .D(n61), .E(n1219), .CK(clk), 
        .Q(n60) );
  EDFFTRX1 index_buffer_reg_14__4_ ( .RN(n1203), .D(n60), .E(n12201), .CK(clk), 
        .Q(n59) );
  EDFFTRX1 index_buffer_reg_13__4_ ( .RN(n1203), .D(n59), .E(n1177), .CK(clk), 
        .Q(n58) );
  EDFFTRX1 index_buffer_reg_12__4_ ( .RN(n1203), .D(n58), .E(n12201), .CK(clk), 
        .Q(n57) );
  EDFFTRX1 index_buffer_reg_11__4_ ( .RN(n1203), .D(n57), .E(n1219), .CK(clk), 
        .Q(n56) );
  EDFFTRX1 index_buffer_reg_10__4_ ( .RN(n1203), .D(n56), .E(n1177), .CK(clk), 
        .Q(n55) );
  EDFFTRX1 index_buffer_reg_9__4_ ( .RN(n1203), .D(n55), .E(n1219), .CK(clk), 
        .Q(n54) );
  EDFFTRX1 index_buffer_reg_8__4_ ( .RN(n1203), .D(n54), .E(n12201), .CK(clk), 
        .Q(n53) );
  EDFFTRX1 index_buffer_reg_7__4_ ( .RN(n1202), .D(n53), .E(n1177), .CK(clk), 
        .Q(n52) );
  EDFFTRX1 index_buffer_reg_6__4_ ( .RN(n1202), .D(n52), .E(n12201), .CK(clk), 
        .Q(n51) );
  EDFFTRX1 index_buffer_reg_5__4_ ( .RN(n1202), .D(n51), .E(n1219), .CK(clk), 
        .Q(n50) );
  EDFFTRX1 index_buffer_reg_4__4_ ( .RN(n1202), .D(n50), .E(n1177), .CK(clk), 
        .Q(n49) );
  EDFFTRX1 index_buffer_reg_3__4_ ( .RN(n1202), .D(n49), .E(n1178), .CK(clk), 
        .Q(n48) );
  EDFFTRX1 index_buffer_reg_2__4_ ( .RN(n1202), .D(n48), .E(n12201), .CK(clk), 
        .Q(n47) );
  EDFFTRX1 index_buffer_reg_1__4_ ( .RN(n1202), .D(n47), .E(n1177), .CK(clk), 
        .Q(n46) );
  EDFFTRX1 index_buffer_reg_18__3_ ( .RN(n1201), .D(n37), .E(n12201), .CK(clk), 
        .Q(n36) );
  EDFFTRX1 index_buffer_reg_17__3_ ( .RN(n1201), .D(n36), .E(n1177), .CK(clk), 
        .Q(n35) );
  EDFFTRX1 index_buffer_reg_16__3_ ( .RN(n1201), .D(n35), .E(n11801), .CK(clk), 
        .Q(n34) );
  EDFFTRX1 index_buffer_reg_15__3_ ( .RN(n1201), .D(n34), .E(cnt[0]), .CK(clk), 
        .Q(n33) );
  EDFFTRX1 index_buffer_reg_14__3_ ( .RN(n1201), .D(n33), .E(n1177), .CK(clk), 
        .Q(n32) );
  EDFFTRX1 index_buffer_reg_13__3_ ( .RN(n1201), .D(n32), .E(n1181), .CK(clk), 
        .Q(n31) );
  EDFFTRX1 index_buffer_reg_12__3_ ( .RN(n1201), .D(n31), .E(n12201), .CK(clk), 
        .Q(n30) );
  EDFFTRX1 index_buffer_reg_11__3_ ( .RN(n1201), .D(n30), .E(n1177), .CK(clk), 
        .Q(n29) );
  EDFFTRX1 index_buffer_reg_10__3_ ( .RN(n1201), .D(n29), .E(n1182), .CK(clk), 
        .Q(n28) );
  EDFFTRX1 index_buffer_reg_9__3_ ( .RN(n1201), .D(n28), .E(n1219), .CK(clk), 
        .Q(n27) );
  EDFFTRX1 index_buffer_reg_8__3_ ( .RN(n1201), .D(n27), .E(n1177), .CK(clk), 
        .Q(n26) );
  EDFFTRX1 index_buffer_reg_1__3_ ( .RN(n1205), .D(n20), .E(n1183), .CK(clk), 
        .Q(n19) );
  DFFTRX1 cnt_reg_0_ ( .D(N114), .RN(n1187), .CK(clk), .Q(cnt[0]), .QN(n314)
         );
  EDFFTRX1 index_buffer_reg_0__1_ ( .RN(n1192), .D(n1810), .E(n1183), .CK(clk), 
        .Q(n1431), .QN(n937) );
  EDFFTRX1 index_buffer_reg_0__6_ ( .RN(n1206), .D(n100), .E(n11801), .CK(clk), 
        .Q(n1427), .QN(n935) );
  EDFFTRX1 index_buffer_reg_0__5_ ( .RN(n1204), .D(n730), .E(n12201), .CK(clk), 
        .Q(n1428), .QN(n931) );
  EDFFTRX1 index_buffer_reg_0__7_ ( .RN(n1196), .D(n127), .E(n1179), .CK(clk), 
        .Q(n1426), .QN(n929) );
  EDFFTRX1 index_buffer_reg_0__0_ ( .RN(n1194), .D(n208), .E(n1182), .CK(clk), 
        .Q(n1432), .QN(n927) );
  EDFFTRX1 index_buffer_reg_0__3_ ( .RN(n11901), .D(n19), .E(n1219), .CK(clk), 
        .Q(n1430), .QN(n925) );
  EDFFTRX1 index_buffer_reg_0__4_ ( .RN(n1202), .D(n46), .E(n1181), .CK(clk), 
        .Q(n1429), .QN(n923) );
  DFFX1 index_buffer_reg_32__7_ ( .D(n779), .CK(clk), .QN(n629) );
  DFFX1 index_buffer_reg_32__6_ ( .D(n7801), .CK(clk), .QN(n630) );
  DFFX1 index_buffer_reg_32__5_ ( .D(n781), .CK(clk), .Q(n1324), .QN(n631) );
  DFFX1 index_buffer_reg_32__4_ ( .D(n782), .CK(clk), .Q(n1323), .QN(n632) );
  DFFX1 index_buffer_reg_32__3_ ( .D(n783), .CK(clk), .Q(n1329), .QN(n633) );
  DFFX1 index_buffer_reg_32__2_ ( .D(n784), .CK(clk), .Q(n1328), .QN(n634) );
  DFFX1 index_buffer_reg_32__1_ ( .D(n785), .CK(clk), .QN(n635) );
  DFFX1 index_buffer_reg_32__0_ ( .D(n786), .CK(clk), .QN(n636) );
  DFFX1 index_buffer_reg_31__7_ ( .D(n771), .CK(clk), .QN(n621) );
  DFFX1 index_buffer_reg_31__6_ ( .D(n772), .CK(clk), .QN(n622) );
  DFFX1 index_buffer_reg_31__5_ ( .D(n773), .CK(clk), .Q(n1344), .QN(n623) );
  DFFX1 index_buffer_reg_31__4_ ( .D(n774), .CK(clk), .Q(n1343), .QN(n624) );
  DFFX1 index_buffer_reg_31__3_ ( .D(n775), .CK(clk), .Q(n1349), .QN(n625) );
  DFFX1 index_buffer_reg_31__2_ ( .D(n776), .CK(clk), .Q(n1348), .QN(n626) );
  DFFX1 index_buffer_reg_31__1_ ( .D(n777), .CK(clk), .QN(n627) );
  DFFX1 index_buffer_reg_31__0_ ( .D(n778), .CK(clk), .QN(n628) );
  DFFX1 index_buffer_reg_30__7_ ( .D(n763), .CK(clk), .QN(n613) );
  DFFX1 index_buffer_reg_30__6_ ( .D(n764), .CK(clk), .QN(n614) );
  DFFX1 index_buffer_reg_30__5_ ( .D(n765), .CK(clk), .Q(n1364), .QN(n615) );
  DFFX1 index_buffer_reg_30__4_ ( .D(n766), .CK(clk), .Q(n1363), .QN(n616) );
  DFFX1 index_buffer_reg_30__3_ ( .D(n767), .CK(clk), .Q(n1369), .QN(n617) );
  DFFX1 index_buffer_reg_30__2_ ( .D(n768), .CK(clk), .Q(n1368), .QN(n618) );
  DFFX1 index_buffer_reg_30__1_ ( .D(n769), .CK(clk), .QN(n619) );
  DFFX1 index_buffer_reg_30__0_ ( .D(n7701), .CK(clk), .QN(n620) );
  DFFTRX1 read_addr_low_reg_4_ ( .D(N153), .RN(n1188), .CK(clk), .Q(
        read_addr_low[4]) );
  DFFTRX1 read_addr_low_reg_3_ ( .D(N152), .RN(n796), .CK(clk), .Q(
        read_addr_low[3]) );
  DFFTRX1 rom_a_low_reg_0_ ( .D(N118), .RN(n796), .CK(clk), .Q(rom_a_low[0])
         );
  DFFX1 rd_buffer_reg_0_ ( .D(n795), .CK(clk), .QN(n1263) );
  DFFX1 re_cs_reg_0_ ( .D(N181), .CK(clk), .Q(re_cs[0]), .QN(n1395) );
  DFFX1 rd_buffer_reg_6_ ( .D(n789), .CK(clk), .Q(rd_buffer[6]), .QN(n1289) );
  DFFX1 rd_buffer_reg_5_ ( .D(n7901), .CK(clk), .Q(rd_buffer[5]), .QN(n1287)
         );
  DFFX1 rd_buffer_reg_4_ ( .D(n791), .CK(clk), .Q(rd_buffer[4]), .QN(n1285) );
  DFFX1 rd_buffer_reg_3_ ( .D(n792), .CK(clk), .Q(rd_buffer[3]), .QN(n1283) );
  DFFX1 rd_buffer_reg_2_ ( .D(n793), .CK(clk), .Q(rd_buffer[2]), .QN(n1280) );
  DFFX1 rd_buffer_reg_1_ ( .D(n794), .CK(clk), .Q(rd_buffer[1]), .QN(n1276) );
  DFFX1 write_addr_low_reg_1_ ( .D(N165), .CK(clk), .Q(write_addr_low[1]), 
        .QN(N150) );
  EDFFTRXL index_buffer_reg_27__7_ ( .RN(n1437), .D(index_buffer_28__7_), .E(
        n1182), .CK(clk), .Q(n1530) );
  EDFFTRXL index_buffer_reg_26__7_ ( .RN(n1437), .D(n1530), .E(n1183), .CK(clk), .Q(n1520) );
  EDFFTRXL index_buffer_reg_25__7_ ( .RN(n1438), .D(n1520), .E(n1178), .CK(clk), .Q(n1510) );
  EDFFTRXL index_buffer_reg_24__7_ ( .RN(n1437), .D(n1510), .E(n1179), .CK(clk), .Q(n1500) );
  EDFFTRXL index_buffer_reg_23__7_ ( .RN(n1437), .D(n1500), .E(n11801), .CK(
        clk), .Q(n1490) );
  EDFFTRXL index_buffer_reg_22__7_ ( .RN(n1438), .D(n1490), .E(n1178), .CK(clk), .Q(n1480) );
  EDFFTRXL index_buffer_reg_21__7_ ( .RN(n1437), .D(n1480), .E(n1179), .CK(clk), .Q(n1470) );
  EDFFTRXL index_buffer_reg_3__2_ ( .RN(n1438), .D(n1570), .E(n1181), .CK(clk), 
        .Q(n1560) );
  EDFFTRXL index_buffer_reg_2__2_ ( .RN(n1437), .D(n1560), .E(n1182), .CK(clk), 
        .Q(n1550) );
  EDFFTRXL index_buffer_reg_1__2_ ( .RN(n1438), .D(n1550), .E(n1183), .CK(clk), 
        .Q(n1540) );
  EDFFTRXL index_buffer_reg_13__2_ ( .RN(n1437), .D(n167), .E(n1183), .CK(clk), 
        .Q(n1660) );
  EDFFTRXL index_buffer_reg_12__2_ ( .RN(n1437), .D(n1660), .E(n1181), .CK(clk), .Q(n1650) );
  EDFFTRXL index_buffer_reg_11__2_ ( .RN(n1438), .D(n1650), .E(n1182), .CK(clk), .Q(n1640) );
  EDFFTRXL index_buffer_reg_10__2_ ( .RN(n1438), .D(n1640), .E(n1183), .CK(clk), .Q(n1630) );
  EDFFTRXL index_buffer_reg_9__2_ ( .RN(n1438), .D(n1630), .E(n1181), .CK(clk), 
        .Q(n1620) );
  EDFFTRXL index_buffer_reg_8__2_ ( .RN(n1437), .D(n1620), .E(n1182), .CK(clk), 
        .Q(n1610) );
  EDFFTRXL index_buffer_reg_7__2_ ( .RN(n1437), .D(n1610), .E(n1183), .CK(clk), 
        .Q(n1600) );
  EDFFTRXL index_buffer_reg_6__2_ ( .RN(n1437), .D(n1600), .E(n1181), .CK(clk), 
        .Q(n159) );
  EDFFTRXL index_buffer_reg_5__2_ ( .RN(n1438), .D(n159), .E(n1182), .CK(clk), 
        .Q(n1580) );
  EDFFTRXL index_buffer_reg_27__6_ ( .RN(n1438), .D(index_buffer_28__6_), .E(
        n11801), .CK(clk), .Q(n126) );
  EDFFTRXL index_buffer_reg_26__6_ ( .RN(n1437), .D(n126), .E(n1178), .CK(clk), 
        .Q(n125) );
  EDFFTRXL index_buffer_reg_25__6_ ( .RN(n1438), .D(n125), .E(n1179), .CK(clk), 
        .Q(n12400) );
  EDFFTRXL index_buffer_reg_24__6_ ( .RN(n1438), .D(n12400), .E(n11801), .CK(
        clk), .Q(n12300) );
  EDFFTRXL index_buffer_reg_23__6_ ( .RN(n1437), .D(n12300), .E(n1178), .CK(
        clk), .Q(n12200) );
  EDFFTRXL index_buffer_reg_22__6_ ( .RN(n1438), .D(n12200), .E(n1179), .CK(
        clk), .Q(n12100) );
  EDFFTRXL index_buffer_reg_21__6_ ( .RN(n1438), .D(n12100), .E(n11801), .CK(
        clk), .Q(n12000) );
  EDFFTRXL index_buffer_reg_20__7_ ( .RN(n1437), .D(n1470), .E(n11801), .CK(
        clk), .Q(n1460) );
  EDFFTRXL index_buffer_reg_20__6_ ( .RN(n1437), .D(n12000), .E(n1178), .CK(
        clk), .Q(n11900) );
  EDFFTRXL index_buffer_reg_19__7_ ( .RN(n1438), .D(n1460), .E(n1178), .CK(clk), .Q(n1450) );
  EDFFTRXL index_buffer_reg_19__6_ ( .RN(n1438), .D(n11900), .E(n1179), .CK(
        clk), .Q(n11800) );
  EDFFTRXL index_buffer_reg_18__7_ ( .RN(n1437), .D(n1450), .E(n1179), .CK(clk), .Q(n1440) );
  EDFFTRXL index_buffer_reg_18__6_ ( .RN(n1438), .D(n11800), .E(n11801), .CK(
        clk), .Q(n1170) );
  EDFFTRXL index_buffer_reg_17__7_ ( .RN(n1437), .D(n1440), .E(n11801), .CK(
        clk), .Q(n14340) );
  EDFFTRXL index_buffer_reg_17__6_ ( .RN(n1437), .D(n1170), .E(n1178), .CK(clk), .Q(n1160) );
  EDFFTRXL index_buffer_reg_16__7_ ( .RN(n1438), .D(n14340), .E(n1178), .CK(
        clk), .Q(n14210) );
  EDFFTRXL index_buffer_reg_16__6_ ( .RN(n1438), .D(n1160), .E(n1179), .CK(clk), .Q(n1150) );
  EDFFTRXL index_buffer_reg_15__7_ ( .RN(n1437), .D(n14210), .E(n1179), .CK(
        clk), .Q(n14100) );
  EDFFTRXL index_buffer_reg_15__6_ ( .RN(n1438), .D(n1150), .E(n11801), .CK(
        clk), .Q(n11400) );
  EDFFTRXL index_buffer_reg_14__7_ ( .RN(n1437), .D(n14100), .E(n11801), .CK(
        clk), .Q(n14000) );
  EDFFTRXL index_buffer_reg_14__6_ ( .RN(n1437), .D(n11400), .E(n1178), .CK(
        clk), .Q(n113) );
  EDFFTRXL index_buffer_reg_13__7_ ( .RN(n1438), .D(n14000), .E(n1178), .CK(
        clk), .Q(n13900) );
  EDFFTRXL index_buffer_reg_13__6_ ( .RN(n1438), .D(n113), .E(n1179), .CK(clk), 
        .Q(n112) );
  EDFFTRXL index_buffer_reg_12__7_ ( .RN(n1438), .D(n13900), .E(n1179), .CK(
        clk), .Q(n13800) );
  EDFFTRXL index_buffer_reg_12__6_ ( .RN(n1437), .D(n112), .E(n11801), .CK(clk), .Q(n111) );
  EDFFTRXL index_buffer_reg_11__7_ ( .RN(n1438), .D(n13800), .E(n11801), .CK(
        clk), .Q(n137) );
  EDFFTRXL index_buffer_reg_11__6_ ( .RN(n1437), .D(n111), .E(n1178), .CK(clk), 
        .Q(n110) );
  EDFFTRXL index_buffer_reg_10__7_ ( .RN(n1438), .D(n137), .E(n1178), .CK(clk), 
        .Q(n136) );
  EDFFTRXL index_buffer_reg_10__6_ ( .RN(n1437), .D(n110), .E(n1179), .CK(clk), 
        .Q(n109) );
  EDFFTRXL index_buffer_reg_9__7_ ( .RN(n1437), .D(n136), .E(n1179), .CK(clk), 
        .Q(n135) );
  EDFFTRXL index_buffer_reg_9__6_ ( .RN(n1438), .D(n109), .E(n11801), .CK(clk), 
        .Q(n108) );
  EDFFTRXL index_buffer_reg_8__7_ ( .RN(n1437), .D(n135), .E(n11801), .CK(clk), 
        .Q(n134) );
  EDFFTRXL index_buffer_reg_8__6_ ( .RN(n1437), .D(n108), .E(n1178), .CK(clk), 
        .Q(n107) );
  EDFFTRXL index_buffer_reg_7__7_ ( .RN(n1438), .D(n134), .E(n1178), .CK(clk), 
        .Q(n133) );
  EDFFTRXL index_buffer_reg_7__6_ ( .RN(n1438), .D(n107), .E(n1179), .CK(clk), 
        .Q(n106) );
  EDFFTRXL index_buffer_reg_6__7_ ( .RN(n1438), .D(n133), .E(n1179), .CK(clk), 
        .Q(n132) );
  EDFFTRXL index_buffer_reg_5__7_ ( .RN(n1437), .D(n132), .E(n11801), .CK(clk), 
        .Q(n131) );
  EDFFTRXL index_buffer_reg_4__7_ ( .RN(n1437), .D(n131), .E(n1178), .CK(clk), 
        .Q(n130) );
  EDFFTRXL index_buffer_reg_3__7_ ( .RN(n1438), .D(n130), .E(n1179), .CK(clk), 
        .Q(n129) );
  EDFFTRXL index_buffer_reg_2__7_ ( .RN(n1437), .D(n129), .E(n11801), .CK(clk), 
        .Q(n128) );
  EDFFTRXL index_buffer_reg_1__7_ ( .RN(n1438), .D(n128), .E(n1178), .CK(clk), 
        .Q(n127) );
  EDFFTRXL rd_buffer_reg_37_ ( .RN(n1437), .D(n239), .E(n1221), .CK(clk), .Q(
        n238) );
  EDFFTRXL rd_buffer_reg_36_ ( .RN(n1438), .D(n240), .E(n1221), .CK(clk), .Q(
        n239) );
  EDFFTRXL rd_buffer_reg_35_ ( .RN(n1437), .D(n241), .E(n1221), .CK(clk), .Q(
        n240) );
  EDFFTRX1 rd_buffer_reg_40_ ( .RN(n1438), .D(rd_buffer[39]), .E(n1221), .CK(
        clk), .Q(rd_buffer[40]), .QN(n1295) );
  DFFX1 index_buffer_reg_29__5_ ( .D(n757), .CK(clk), .QN(n1236) );
  DFFX1 index_buffer_reg_29__3_ ( .D(n759), .CK(clk), .QN(n1239) );
  DFFX1 index_buffer_reg_29__1_ ( .D(n761), .CK(clk), .QN(n12401) );
  DFFX1 index_buffer_reg_28__6_ ( .D(n748), .CK(clk), .Q(index_buffer_28__6_), 
        .QN(n1237) );
  DFFX1 index_buffer_reg_29__7_ ( .D(n755), .CK(clk), .QN(n1238) );
  DFFX1 index_buffer_reg_28__5_ ( .D(n749), .CK(clk), .Q(index_buffer_28__5_), 
        .QN(n599) );
  DFFX1 index_buffer_reg_28__3_ ( .D(n751), .CK(clk), .Q(index_buffer_28__3_), 
        .QN(n601) );
  DFFTRX1 rw_reg ( .D(N138), .RN(n1187), .CK(clk), .Q(rw), .QN(n1433) );
  DFFTRX1 write_addr_low_reg_3_ ( .D(N142), .RN(n1188), .CK(clk), .Q(
        write_addr_low[3]), .QN(n1243) );
  XOR2X1 U223 ( .A(n1257), .B(write_addr_high[3]), .Y(n1253) );
  XOR2X1 U224 ( .A(n1257), .B(write_addr_high[4]), .Y(n1249) );
  OAI222XL U225 ( .A0(n1296), .A1(n1304), .B0(n366), .B1(n1298), .C0(n630), 
        .C1(n1185), .Y(n7801) );
  OAI222XL U226 ( .A0(n1296), .A1(n1305), .B0(n365), .B1(n1298), .C0(n629), 
        .C1(n1186), .Y(n779) );
  NOR2X2 U227 ( .A(n1184), .B(n802), .Y(n796) );
  OA21XL U228 ( .A0(n1433), .A1(n1255), .B0(n1256), .Y(n797) );
  OA21XL U229 ( .A0(sram_wen), .A1(n1249), .B0(n1250), .Y(n798) );
  OA21XL U230 ( .A0(n828), .A1(n1253), .B0(n1254), .Y(n799) );
  AOI21X1 U231 ( .A0(rw), .A1(n944), .B0(n1141), .Y(n8001) );
  INVX1 U232 ( .A(reset), .Y(n801) );
  INVX3 U233 ( .A(n801), .Y(n802) );
  XOR2X1 U235 ( .A(n1257), .B(write_addr_high[2]), .Y(n1255) );
  OAI222XL U236 ( .A0(index_buffer_28__5_), .A1(n1236), .B0(
        index_buffer_28__5_), .B1(n1222), .C0(n1236), .C1(n1222), .Y(n1223) );
  OA22XL U237 ( .A0(n1224), .A1(index_buffer_28__3_), .B0(n1224), .B1(n1239), 
        .Y(n1228) );
  INVXL U238 ( .A(n1307), .Y(n807) );
  INVX3 U239 ( .A(n807), .Y(n808) );
  INVXL U240 ( .A(n1333), .Y(n809) );
  INVX3 U241 ( .A(n809), .Y(n8101) );
  INVXL U242 ( .A(n1353), .Y(n811) );
  INVX3 U243 ( .A(n811), .Y(n812) );
  INVXL U244 ( .A(n1420), .Y(n813) );
  INVX12 U245 ( .A(n813), .Y(sram_a[6]) );
  OAI2BB1X1 U246 ( .A0N(rw), .A1N(n943), .B0(n1142), .Y(n1420) );
  INVXL U247 ( .A(n1423), .Y(n815) );
  INVX12 U248 ( .A(n815), .Y(sram_a[2]) );
  OAI2BB1X1 U249 ( .A0N(rw), .A1N(n946), .B0(n1138), .Y(n1423) );
  INVX12 U250 ( .A(n8001), .Y(sram_a[5]) );
  INVXL U251 ( .A(n1424), .Y(n818) );
  INVX12 U252 ( .A(n818), .Y(sram_a[1]) );
  OAI2BB1X1 U253 ( .A0N(rw), .A1N(n945), .B0(n1137), .Y(n1424) );
  INVX12 U254 ( .A(n798), .Y(sram_a[9]) );
  INVXL U255 ( .A(n1425), .Y(n821) );
  INVX12 U256 ( .A(n821), .Y(sram_a[0]) );
  AO21X1 U257 ( .A0(rw), .A1(n947), .B0(n11401), .Y(n1425) );
  INVX12 U258 ( .A(n799), .Y(sram_a[8]) );
  INVX12 U259 ( .A(n797), .Y(sram_a[7]) );
  CLKINVX1 U261 ( .A(n1433), .Y(n826) );
  INVX12 U262 ( .A(n826), .Y(sram_wen) );
  CLKINVX2 U263 ( .A(n826), .Y(n828) );
  BUFX12 U265 ( .A(n1417), .Y(rom_a[2]) );
  BUFX12 U266 ( .A(n1416), .Y(rom_a[3]) );
  XOR2XL U267 ( .A(rom_a_high[1]), .B(re_cs[2]), .Y(n1416) );
  BUFX12 U268 ( .A(n1415), .Y(rom_a[4]) );
  XOR2XL U269 ( .A(rom_a_high[2]), .B(re_cs[2]), .Y(n1415) );
  BUFX12 U270 ( .A(n1414), .Y(rom_a[5]) );
  XOR2XL U271 ( .A(rom_a_high[3]), .B(re_cs[2]), .Y(n1414) );
  BUFX12 U272 ( .A(n1413), .Y(rom_a[6]) );
  XOR2XL U273 ( .A(rom_a_high[4]), .B(re_cs[2]), .Y(n1413) );
  BUFX12 U274 ( .A(n1422), .Y(sram_a[3]) );
  BUFX12 U275 ( .A(n1421), .Y(sram_a[4]) );
  NAND2X2 U276 ( .A(n1314), .B(n1335), .Y(n1332) );
  NAND2X2 U277 ( .A(n1314), .B(n1355), .Y(n1352) );
  NAND2X2 U278 ( .A(n1314), .B(n1315), .Y(n1306) );
  XNOR2X1 U279 ( .A(n1257), .B(write_addr_high[1]), .Y(n943) );
  OAI2BB1X2 U280 ( .A0N(N397), .A1N(rd_buffer[12]), .B0(n1292), .Y(n1373) );
  XNOR2X1 U281 ( .A(n942), .B(write_addr_low[2]), .Y(n946) );
  XNOR2X1 U282 ( .A(n1242), .B(re_cs[2]), .Y(n944) );
  INVX12 U283 ( .A(n923), .Y(sram_d[4]) );
  OAI222XL U284 ( .A0(n1296), .A1(n1300), .B0(n370), .B1(n1298), .C0(n634), 
        .C1(n1185), .Y(n784) );
  OAI222XL U285 ( .A0(n1296), .A1(n1301), .B0(n369), .B1(n1298), .C0(n633), 
        .C1(n1185), .Y(n783) );
  OAI222XL U286 ( .A0(n1296), .A1(n1302), .B0(n368), .B1(n1298), .C0(n632), 
        .C1(n1186), .Y(n782) );
  OAI222XL U287 ( .A0(n1296), .A1(n1303), .B0(n367), .B1(n1298), .C0(n631), 
        .C1(n1185), .Y(n781) );
  NAND3X2 U288 ( .A(rd_buffer[7]), .B(n1292), .C(rd_sram), .Y(n1296) );
  XNOR2X1 U289 ( .A(n942), .B(write_addr_low[1]), .Y(n945) );
  INVX12 U290 ( .A(n925), .Y(sram_d[3]) );
  INVX12 U291 ( .A(n927), .Y(sram_d[0]) );
  INVX12 U292 ( .A(n929), .Y(sram_d[7]) );
  XNOR2X1 U293 ( .A(n942), .B(N149), .Y(n947) );
  NAND3BX2 U294 ( .AN(rd_sram), .B(n1292), .C(rd_buffer[7]), .Y(n1298) );
  AOI31X4 U295 ( .A0(rd_buffer[12]), .A1(n11901), .A2(N397), .B0(n1144), .Y(
        n1372) );
  INVX12 U296 ( .A(n931), .Y(sram_d[5]) );
  NAND4X1 U297 ( .A(n1175), .B(n1134), .C(n1135), .D(n1136), .Y(n933) );
  INVX12 U298 ( .A(n933), .Y(finish) );
  INVX12 U299 ( .A(n935), .Y(sram_d[6]) );
  INVX12 U300 ( .A(n937), .Y(sram_d[1]) );
  BUFX12 U301 ( .A(n1418), .Y(rom_a[1]) );
  XOR2XL U302 ( .A(rom_a_low[1]), .B(n941), .Y(n1418) );
  BUFX12 U303 ( .A(n1419), .Y(rom_a[0]) );
  XOR2XL U304 ( .A(rom_a_low[0]), .B(n941), .Y(n1419) );
  INVX1 U305 ( .A(n1429), .Y(n1310) );
  INVX1 U306 ( .A(n1428), .Y(n1311) );
  NOR2XL U307 ( .A(n1431), .B(n635), .Y(n1331) );
  AOI211XL U308 ( .A0(n1431), .A1(n635), .B0(n1432), .C0(n636), .Y(n1330) );
  NOR2XL U309 ( .A(n1431), .B(n619), .Y(n1371) );
  AOI211XL U310 ( .A0(n619), .A1(n1431), .B0(n1432), .C0(n620), .Y(n1370) );
  NOR2XL U311 ( .A(n1431), .B(n627), .Y(n1351) );
  AOI211XL U312 ( .A0(n627), .A1(n1431), .B0(n1432), .C0(n628), .Y(n1350) );
  NAND2XL U313 ( .A(n1428), .B(n631), .Y(n1318) );
  NAND2XL U314 ( .A(n615), .B(n1428), .Y(n1358) );
  NAND2XL U315 ( .A(n623), .B(n1428), .Y(n1338) );
  AO21XL U316 ( .A0(n613), .A1(n1426), .B0(n1356), .Y(n1354) );
  AOI22XL U317 ( .A0(n614), .A1(n1427), .B0(n616), .B1(n1429), .Y(n1359) );
  AO21XL U318 ( .A0(n621), .A1(n1426), .B0(n1336), .Y(n1334) );
  AOI22XL U319 ( .A0(n622), .A1(n1427), .B0(n624), .B1(n1429), .Y(n1339) );
  AO21XL U320 ( .A0(n1426), .A1(n629), .B0(n1316), .Y(n1313) );
  AOI22XL U321 ( .A0(n1427), .A1(n630), .B0(n1429), .B1(n632), .Y(n1319) );
  NAND4XL U322 ( .A(n947), .B(n945), .C(n1404), .D(n946), .Y(n1403) );
  NOR2XL U323 ( .A(n1258), .B(n1261), .Y(n1404) );
  NAND3XL U324 ( .A(n1261), .B(n1258), .C(n1407), .Y(n14001) );
  NOR3XL U325 ( .A(n946), .B(n945), .C(n947), .Y(n1407) );
  NOR3XL U326 ( .A(n942), .B(n1257), .C(n1395), .Y(n13901) );
  INVX3 U327 ( .A(n1176), .Y(n1177) );
  NAND4XL U328 ( .A(n1255), .B(n1253), .C(n1249), .D(n1405), .Y(n1401) );
  NOR3XL U329 ( .A(n943), .B(n828), .C(n944), .Y(n1405) );
  NAND4BXL U330 ( .AN(n1255), .B(n943), .C(n944), .D(n1406), .Y(n1402) );
  NOR3XL U331 ( .A(n1253), .B(n828), .C(n1249), .Y(n1406) );
  CLKINVX1 U332 ( .A(n1219), .Y(n1176) );
  AND2XL U333 ( .A(add_95_carry[4]), .B(write_addr_low[4]), .Y(add_95_carry[5]) );
  AND2XL U334 ( .A(write_addr_low[1]), .B(write_addr_low[2]), .Y(
        add_95_carry[3]) );
  AND2XL U335 ( .A(add_95_carry[6]), .B(write_addr_high[1]), .Y(
        add_95_carry[7]) );
  XOR2XL U336 ( .A(write_addr_low[4]), .B(add_95_carry[4]), .Y(N153) );
  XOR2XL U337 ( .A(write_addr_high[1]), .B(add_95_carry[6]), .Y(N155) );
  XOR2XL U338 ( .A(write_addr_low[2]), .B(write_addr_low[1]), .Y(N151) );
  CLKBUFX3 U339 ( .A(n1209), .Y(n1201) );
  CLKBUFX3 U340 ( .A(n1209), .Y(n1202) );
  CLKBUFX3 U341 ( .A(n1208), .Y(n1203) );
  CLKBUFX3 U342 ( .A(n1208), .Y(n1204) );
  CLKBUFX3 U343 ( .A(n1207), .Y(n1205) );
  CLKBUFX3 U344 ( .A(n1207), .Y(n1206) );
  CLKBUFX3 U346 ( .A(n1213), .Y(n1192) );
  CLKBUFX3 U348 ( .A(n1213), .Y(n1194) );
  CLKBUFX3 U350 ( .A(n1212), .Y(n1196) );
  CLKBUFX3 U352 ( .A(n1211), .Y(n1198) );
  CLKBUFX3 U353 ( .A(n12101), .Y(n1199) );
  CLKBUFX3 U354 ( .A(n12101), .Y(n12001) );
  CLKBUFX3 U355 ( .A(n1214), .Y(n11901) );
  CLKBUFX3 U356 ( .A(n1215), .Y(n1214) );
  CLKBUFX3 U357 ( .A(n1217), .Y(n1209) );
  CLKBUFX3 U358 ( .A(n1217), .Y(n1208) );
  CLKBUFX3 U359 ( .A(n1217), .Y(n1207) );
  CLKBUFX3 U360 ( .A(n1215), .Y(n1213) );
  CLKBUFX3 U361 ( .A(n1216), .Y(n1212) );
  CLKBUFX3 U362 ( .A(n1216), .Y(n1211) );
  CLKBUFX3 U363 ( .A(n1216), .Y(n12101) );
  CLKBUFX3 U364 ( .A(n796), .Y(n1188) );
  CLKBUFX3 U365 ( .A(n1218), .Y(n1215) );
  INVX3 U366 ( .A(n1144), .Y(n1185) );
  INVX3 U367 ( .A(n1144), .Y(n1186) );
  CLKBUFX3 U368 ( .A(n1216), .Y(n1217) );
  CLKBUFX3 U369 ( .A(n1218), .Y(n1216) );
  BUFX4 U370 ( .A(n1411), .Y(n1184) );
  CLKINVX1 U371 ( .A(n1397), .Y(n1411) );
  CLKBUFX3 U372 ( .A(n796), .Y(n1187) );
  CLKBUFX3 U373 ( .A(n1437), .Y(n1218) );
  INVX4 U374 ( .A(n314), .Y(n11801) );
  INVX4 U375 ( .A(n314), .Y(n1179) );
  INVX4 U376 ( .A(n1176), .Y(n1178) );
  INVX4 U377 ( .A(n314), .Y(n1183) );
  INVX4 U378 ( .A(n1176), .Y(n1182) );
  INVX4 U379 ( .A(n1176), .Y(n1181) );
  AND4X1 U380 ( .A(n1246), .B(n1245), .C(n1374), .D(n1244), .Y(n1134) );
  AND3X2 U381 ( .A(n1248), .B(n1247), .C(times[0]), .Y(n1135) );
  AND2X2 U382 ( .A(times[2]), .B(times[1]), .Y(n1136) );
  AND4X1 U383 ( .A(n1375), .B(n1376), .C(n1377), .D(n1378), .Y(n1175) );
  MXI2X1 U384 ( .A(n1259), .B(n1260), .S0(read_addr_low[1]), .Y(n1137) );
  MXI2X1 U385 ( .A(n1259), .B(n1260), .S0(read_addr_low[2]), .Y(n1138) );
  OAI21XL U386 ( .A0(n828), .A1(n1261), .B0(n1139), .Y(n1422) );
  MXI2X1 U387 ( .A(n1259), .B(n1260), .S0(read_addr_low[3]), .Y(n1139) );
  CLKMX2X2 U388 ( .A(n1259), .B(n1260), .S0(read_addr_low[0]), .Y(n11401) );
  CLKMX2X2 U389 ( .A(n1251), .B(n1252), .S0(read_addr_high[0]), .Y(n1141) );
  MXI2X1 U390 ( .A(n1251), .B(n1252), .S0(read_addr_high[1]), .Y(n1142) );
  OAI21XL U391 ( .A0(n828), .A1(n1258), .B0(n1143), .Y(n1421) );
  MXI2X1 U392 ( .A(n1259), .B(n1260), .S0(read_addr_low[4]), .Y(n1143) );
  CLKINVX2 U393 ( .A(n1430), .Y(n1309) );
  NOR2X2 U394 ( .A(n802), .B(n1144), .Y(n1292) );
  AND2X2 U395 ( .A(n314), .B(n11901), .Y(n1144) );
  CLKBUFX3 U396 ( .A(cnt[0]), .Y(n1219) );
  CLKBUFX8 U397 ( .A(cnt[0]), .Y(n1221) );
  CLKBUFX3 U398 ( .A(cnt[0]), .Y(n12201) );
  XOR2X1 U399 ( .A(write_addr_high[4]), .B(add_95_carry[9]), .Y(N158) );
  AND2X1 U400 ( .A(add_95_carry[8]), .B(write_addr_high[3]), .Y(
        add_95_carry[9]) );
  XOR2X1 U401 ( .A(write_addr_high[3]), .B(add_95_carry[8]), .Y(N157) );
  AND2X1 U402 ( .A(add_95_carry[7]), .B(write_addr_high[2]), .Y(
        add_95_carry[8]) );
  XOR2X1 U403 ( .A(write_addr_high[2]), .B(add_95_carry[7]), .Y(N156) );
  OR2X1 U404 ( .A(write_addr_high[0]), .B(add_95_carry[5]), .Y(add_95_carry[6]) );
  XNOR2X1 U405 ( .A(add_95_carry[5]), .B(write_addr_high[0]), .Y(N154) );
  AND2X1 U406 ( .A(add_95_carry[3]), .B(write_addr_low[3]), .Y(add_95_carry[4]) );
  XOR2X1 U407 ( .A(write_addr_low[3]), .B(add_95_carry[3]), .Y(N152) );
  NAND2BX1 U408 ( .AN(index_buffer_28__4_), .B(index_buffer_29__4_), .Y(n1222)
         );
  OAI222XL U409 ( .A0(index_buffer_29__6_), .A1(n1223), .B0(n1237), .B1(n1223), 
        .C0(index_buffer_29__6_), .C1(n1237), .Y(n1234) );
  NAND2BX1 U410 ( .AN(index_buffer_28__2_), .B(index_buffer_29__2_), .Y(n1226)
         );
  OAI22XL U411 ( .A0(index_buffer_28__3_), .A1(n1239), .B0(index_buffer_28__3_), .B1(n1226), .Y(n1232) );
  NOR2BX1 U412 ( .AN(index_buffer_28__2_), .B(index_buffer_29__2_), .Y(n1224)
         );
  AOI21X1 U413 ( .A0(index_buffer_28__1_), .A1(n12401), .B0(
        index_buffer_28__0_), .Y(n1225) );
  AOI2BB2X1 U414 ( .B0(n1225), .B1(index_buffer_29__0_), .A0N(
        index_buffer_28__1_), .A1N(n12401), .Y(n1227) );
  OAI22XL U415 ( .A0(n1228), .A1(n1227), .B0(n1226), .B1(n1239), .Y(n1231) );
  NOR2BX1 U416 ( .AN(index_buffer_28__4_), .B(index_buffer_29__4_), .Y(n1229)
         );
  OAI22XL U417 ( .A0(n1229), .A1(n1236), .B0(index_buffer_28__5_), .B1(n1229), 
        .Y(n12301) );
  OAI221XL U418 ( .A0(index_buffer_29__6_), .A1(n1237), .B0(n1232), .B1(n1231), 
        .C0(n12301), .Y(n1233) );
  AO22X1 U419 ( .A0(n1238), .A1(index_buffer_28__7_), .B0(n1234), .B1(n1233), 
        .Y(n1235) );
  OAI21XL U420 ( .A0(index_buffer_28__7_), .A1(n1238), .B0(n1235), .Y(N397) );
  MXI2X1 U421 ( .A(n1251), .B(n1252), .S0(read_addr_high[4]), .Y(n1250) );
  MXI2X1 U422 ( .A(n1251), .B(n1252), .S0(read_addr_high[3]), .Y(n1254) );
  MXI2X1 U423 ( .A(n1251), .B(n1252), .S0(read_addr_high[2]), .Y(n1256) );
  NOR2BX1 U424 ( .AN(n828), .B(re_cs[2]), .Y(n1252) );
  NOR2BX1 U425 ( .AN(n828), .B(n1257), .Y(n1251) );
  NOR2BX1 U426 ( .AN(n828), .B(n941), .Y(n1260) );
  NOR2BX1 U427 ( .AN(n828), .B(n942), .Y(n1259) );
  XOR2X1 U428 ( .A(rom_a_high[0]), .B(re_cs[2]), .Y(n1417) );
  MXI2X1 U429 ( .A(n1262), .B(n1263), .S0(n1264), .Y(n795) );
  AOI2BB1X1 U430 ( .A0N(n314), .A1N(n1265), .B0(n802), .Y(n1264) );
  NAND2X1 U431 ( .A(n1266), .B(n11901), .Y(n1262) );
  MXI2X1 U432 ( .A(n1267), .B(n1268), .S0(n941), .Y(n1266) );
  OAI221XL U433 ( .A0(n1269), .A1(n1270), .B0(n1263), .B1(n1271), .C0(n1272), 
        .Y(n794) );
  AOI2BB2X1 U434 ( .B0(rd_buffer[1]), .B1(n1144), .A0N(n1273), .A1N(n1274), 
        .Y(n1272) );
  OAI221XL U435 ( .A0(n1269), .A1(n1275), .B0(n1271), .B1(n1276), .C0(n1277), 
        .Y(n793) );
  AOI2BB2X1 U436 ( .B0(rd_buffer[2]), .B1(n1144), .A0N(n1273), .A1N(n1278), 
        .Y(n1277) );
  OAI221XL U437 ( .A0(n1269), .A1(n1279), .B0(n1271), .B1(n1280), .C0(n1281), 
        .Y(n792) );
  AOI2BB2X1 U438 ( .B0(rd_buffer[3]), .B1(n1144), .A0N(n1273), .A1N(n1282), 
        .Y(n1281) );
  OAI221XL U439 ( .A0(n1269), .A1(n1282), .B0(n1271), .B1(n1283), .C0(n1284), 
        .Y(n791) );
  AOI2BB2X1 U440 ( .B0(rd_buffer[4]), .B1(n1144), .A0N(n1273), .A1N(n1279), 
        .Y(n1284) );
  CLKINVX1 U441 ( .A(rom_q[3]), .Y(n1279) );
  CLKINVX1 U442 ( .A(rom_q[4]), .Y(n1282) );
  OAI221XL U443 ( .A0(n1269), .A1(n1278), .B0(n1271), .B1(n1285), .C0(n1286), 
        .Y(n7901) );
  AOI2BB2X1 U444 ( .B0(rd_buffer[5]), .B1(n1144), .A0N(n1273), .A1N(n1275), 
        .Y(n1286) );
  CLKINVX1 U445 ( .A(rom_q[2]), .Y(n1275) );
  CLKINVX1 U446 ( .A(rom_q[5]), .Y(n1278) );
  OAI221XL U447 ( .A0(n1269), .A1(n1274), .B0(n1271), .B1(n1287), .C0(n1288), 
        .Y(n789) );
  AOI2BB2X1 U448 ( .B0(rd_buffer[6]), .B1(n1144), .A0N(n1270), .A1N(n1273), 
        .Y(n1288) );
  CLKINVX1 U449 ( .A(rom_q[1]), .Y(n1270) );
  CLKINVX1 U450 ( .A(rom_q[6]), .Y(n1274) );
  OAI221XL U451 ( .A0(n1269), .A1(n1268), .B0(n1271), .B1(n1289), .C0(n1290), 
        .Y(n788) );
  AOI2BB2X1 U452 ( .B0(rd_buffer[7]), .B1(n1144), .A0N(n1273), .A1N(n1267), 
        .Y(n1290) );
  CLKINVX1 U453 ( .A(rom_q[0]), .Y(n1267) );
  NAND3X1 U454 ( .A(n1291), .B(n941), .C(n1292), .Y(n1273) );
  NAND2X1 U455 ( .A(n1292), .B(n1265), .Y(n1271) );
  CLKINVX1 U456 ( .A(rom_q[7]), .Y(n1268) );
  NAND3X1 U457 ( .A(n1291), .B(n942), .C(n1292), .Y(n1269) );
  CLKINVX1 U458 ( .A(n1265), .Y(n1291) );
  NAND3X1 U459 ( .A(cnt[2]), .B(cnt[1]), .C(cnt[3]), .Y(n1265) );
  AOI2BB1X1 U460 ( .A0N(n1293), .A1N(n1294), .B0(n802), .Y(n787) );
  NAND3X1 U461 ( .A(rd_buffer[7]), .B(cs), .C(n326), .Y(n1294) );
  NAND3X1 U462 ( .A(n1295), .B(n1408), .C(n1409), .Y(n1293) );
  OAI222XL U463 ( .A0(n1296), .A1(n1297), .B0(n372), .B1(n1298), .C0(n636), 
        .C1(n1186), .Y(n786) );
  CLKINVX1 U464 ( .A(sram_q[0]), .Y(n1297) );
  OAI222XL U465 ( .A0(n1296), .A1(n1299), .B0(n371), .B1(n1298), .C0(n635), 
        .C1(n1186), .Y(n785) );
  CLKINVX1 U466 ( .A(sram_q[1]), .Y(n1299) );
  CLKINVX1 U467 ( .A(sram_q[2]), .Y(n1300) );
  CLKINVX1 U468 ( .A(sram_q[3]), .Y(n1301) );
  CLKINVX1 U469 ( .A(sram_q[4]), .Y(n1302) );
  CLKINVX1 U470 ( .A(sram_q[5]), .Y(n1303) );
  CLKINVX1 U471 ( .A(sram_q[6]), .Y(n1304) );
  CLKINVX1 U472 ( .A(sram_q[7]), .Y(n1305) );
  OAI222XL U473 ( .A0(n1306), .A1(n927), .B0(n636), .B1(n808), .C0(n628), .C1(
        n1186), .Y(n778) );
  OAI222XL U474 ( .A0(n937), .A1(n1306), .B0(n635), .B1(n808), .C0(n627), .C1(
        n1186), .Y(n777) );
  OAI222XL U475 ( .A0(n1308), .A1(n1306), .B0(n634), .B1(n808), .C0(n626), 
        .C1(n1186), .Y(n776) );
  OAI222XL U476 ( .A0(n1309), .A1(n1306), .B0(n633), .B1(n808), .C0(n625), 
        .C1(n1186), .Y(n775) );
  OAI222XL U477 ( .A0(n1310), .A1(n1306), .B0(n632), .B1(n808), .C0(n624), 
        .C1(n1186), .Y(n774) );
  OAI222XL U478 ( .A0(n1311), .A1(n1306), .B0(n631), .B1(n808), .C0(n623), 
        .C1(n1186), .Y(n773) );
  OAI222XL U479 ( .A0(n935), .A1(n1306), .B0(n630), .B1(n808), .C0(n622), .C1(
        n1186), .Y(n772) );
  OAI222XL U480 ( .A0(n929), .A1(n1306), .B0(n629), .B1(n808), .C0(n621), .C1(
        n1186), .Y(n771) );
  OAI221XL U481 ( .A0(n629), .A1(n1312), .B0(n1295), .B1(n1313), .C0(n1292), 
        .Y(n1307) );
  OAI21XL U482 ( .A0(n629), .A1(n1426), .B0(n1313), .Y(n1315) );
  AOI32X1 U483 ( .A0(n1317), .A1(n1318), .A2(n1319), .B0(n1320), .B1(n1321), 
        .Y(n1316) );
  OAI21XL U484 ( .A0(n1322), .A1(n630), .B0(n1427), .Y(n1321) );
  NAND2X1 U485 ( .A(n1322), .B(n630), .Y(n1320) );
  AOI32X1 U486 ( .A0(n1318), .A1(n1310), .A2(n1323), .B0(n1311), .B1(n1324), 
        .Y(n1322) );
  OAI211X1 U487 ( .A0(n633), .A1(n1325), .B0(n1326), .C0(n1327), .Y(n1317) );
  OAI2BB1X1 U488 ( .A0N(n1325), .A1N(n633), .B0(n1309), .Y(n1327) );
  OAI222XL U489 ( .A0(n1328), .A1(n1308), .B0(n1329), .B1(n1309), .C0(n1330), 
        .C1(n1331), .Y(n1326) );
  NAND2X1 U490 ( .A(n1308), .B(n1328), .Y(n1325) );
  OAI222XL U491 ( .A0(n927), .A1(n1332), .B0(n628), .B1(n8101), .C0(n620), 
        .C1(n1186), .Y(n7701) );
  OAI222XL U492 ( .A0(n937), .A1(n1332), .B0(n627), .B1(n8101), .C0(n619), 
        .C1(n1186), .Y(n769) );
  OAI222XL U493 ( .A0(n1308), .A1(n1332), .B0(n626), .B1(n8101), .C0(n618), 
        .C1(n1186), .Y(n768) );
  OAI222XL U494 ( .A0(n1309), .A1(n1332), .B0(n625), .B1(n8101), .C0(n617), 
        .C1(n1186), .Y(n767) );
  OAI222XL U495 ( .A0(n1310), .A1(n1332), .B0(n624), .B1(n8101), .C0(n616), 
        .C1(n1185), .Y(n766) );
  OAI222XL U496 ( .A0(n1311), .A1(n1332), .B0(n623), .B1(n8101), .C0(n615), 
        .C1(n1185), .Y(n765) );
  OAI222XL U497 ( .A0(n935), .A1(n1332), .B0(n622), .B1(n8101), .C0(n614), 
        .C1(n1185), .Y(n764) );
  OAI222XL U498 ( .A0(n929), .A1(n1332), .B0(n621), .B1(n8101), .C0(n613), 
        .C1(n1185), .Y(n763) );
  OAI221XL U499 ( .A0(n621), .A1(n1312), .B0(n1295), .B1(n1334), .C0(n1292), 
        .Y(n1333) );
  OAI21XL U500 ( .A0(n621), .A1(n1426), .B0(n1334), .Y(n1335) );
  AOI32X1 U501 ( .A0(n1337), .A1(n1338), .A2(n1339), .B0(n1340), .B1(n1341), 
        .Y(n1336) );
  OAI21XL U502 ( .A0(n1342), .A1(n622), .B0(n1427), .Y(n1341) );
  NAND2X1 U503 ( .A(n1342), .B(n622), .Y(n1340) );
  AOI32X1 U504 ( .A0(n1338), .A1(n1310), .A2(n1343), .B0(n1311), .B1(n1344), 
        .Y(n1342) );
  OAI211X1 U505 ( .A0(n625), .A1(n1345), .B0(n1346), .C0(n1347), .Y(n1337) );
  OAI2BB1X1 U506 ( .A0N(n1345), .A1N(n625), .B0(n1309), .Y(n1347) );
  OAI222XL U507 ( .A0(n1308), .A1(n1348), .B0(n1309), .B1(n1349), .C0(n1350), 
        .C1(n1351), .Y(n1346) );
  NAND2X1 U508 ( .A(n1308), .B(n1348), .Y(n1345) );
  OAI222XL U509 ( .A0(n927), .A1(n1352), .B0(n620), .B1(n812), .C0(n612), .C1(
        n1185), .Y(n762) );
  OAI222XL U510 ( .A0(n937), .A1(n1352), .B0(n619), .B1(n812), .C0(n12401), 
        .C1(n1185), .Y(n761) );
  OAI222XL U511 ( .A0(n1308), .A1(n1352), .B0(n618), .B1(n812), .C0(n610), 
        .C1(n1185), .Y(n7601) );
  OAI222XL U512 ( .A0(n1309), .A1(n1352), .B0(n617), .B1(n812), .C0(n1239), 
        .C1(n1185), .Y(n759) );
  OAI222XL U513 ( .A0(n1310), .A1(n1352), .B0(n616), .B1(n812), .C0(n608), 
        .C1(n1185), .Y(n758) );
  OAI222XL U514 ( .A0(n1311), .A1(n1352), .B0(n615), .B1(n812), .C0(n1236), 
        .C1(n1185), .Y(n757) );
  OAI222XL U515 ( .A0(n935), .A1(n1352), .B0(n614), .B1(n812), .C0(n606), .C1(
        n1185), .Y(n756) );
  OAI222XL U516 ( .A0(n929), .A1(n1352), .B0(n613), .B1(n812), .C0(n1238), 
        .C1(n1185), .Y(n755) );
  OAI221XL U517 ( .A0(n613), .A1(n1312), .B0(n1295), .B1(n1354), .C0(n1292), 
        .Y(n1353) );
  NAND2X1 U518 ( .A(rd_buffer[40]), .B(n929), .Y(n1312) );
  OAI21XL U519 ( .A0(n613), .A1(n1426), .B0(n1354), .Y(n1355) );
  AOI32X1 U520 ( .A0(n1357), .A1(n1358), .A2(n1359), .B0(n1360), .B1(n1361), 
        .Y(n1356) );
  OAI21XL U521 ( .A0(n1362), .A1(n614), .B0(n1427), .Y(n1361) );
  NAND2X1 U522 ( .A(n1362), .B(n614), .Y(n1360) );
  AOI32X1 U523 ( .A0(n1358), .A1(n1310), .A2(n1363), .B0(n1311), .B1(n1364), 
        .Y(n1362) );
  OAI211X1 U524 ( .A0(n617), .A1(n1365), .B0(n1366), .C0(n1367), .Y(n1357) );
  OAI2BB1X1 U525 ( .A0N(n1365), .A1N(n617), .B0(n1309), .Y(n1367) );
  OAI222XL U526 ( .A0(n1308), .A1(n1368), .B0(n1309), .B1(n1369), .C0(n1370), 
        .C1(n1371), .Y(n1366) );
  NAND2X1 U527 ( .A(n1308), .B(n1368), .Y(n1365) );
  NOR2BX1 U528 ( .AN(n1292), .B(n1295), .Y(n1314) );
  OAI22XL U529 ( .A0(n604), .A1(n1372), .B0(n612), .B1(n1373), .Y(n754) );
  OAI22XL U530 ( .A0(n603), .A1(n1372), .B0(n12401), .B1(n1373), .Y(n753) );
  OAI22XL U531 ( .A0(n602), .A1(n1372), .B0(n610), .B1(n1373), .Y(n752) );
  OAI22XL U532 ( .A0(n601), .A1(n1372), .B0(n1239), .B1(n1373), .Y(n751) );
  OAI22XL U533 ( .A0(n600), .A1(n1372), .B0(n608), .B1(n1373), .Y(n7501) );
  OAI22XL U534 ( .A0(n599), .A1(n1372), .B0(n1236), .B1(n1373), .Y(n749) );
  OAI22XL U535 ( .A0(n1237), .A1(n1372), .B0(n606), .B1(n1373), .Y(n748) );
  OAI22XL U536 ( .A0(n597), .A1(n1372), .B0(n1238), .B1(n1373), .Y(n747) );
  NOR2X1 U538 ( .A(times[16]), .B(times[15]), .Y(n1374) );
  NOR3X1 U539 ( .A(times[7]), .B(times[9]), .C(times[8]), .Y(n1378) );
  NOR3X1 U540 ( .A(times[4]), .B(times[6]), .C(times[5]), .Y(n1377) );
  NOR3X1 U541 ( .A(times[19]), .B(times[3]), .C(times[20]), .Y(n1376) );
  NOR2X1 U542 ( .A(times[18]), .B(times[17]), .Y(n1375) );
  AOI2BB1X1 U543 ( .A0N(n1379), .A1N(n13801), .B0(n802), .Y(N183) );
  OAI21XL U544 ( .A0(n941), .A1(n1257), .B0(n1381), .Y(n13801) );
  OAI2BB1X1 U545 ( .A0N(n1382), .A1N(n1383), .B0(n1384), .Y(n1379) );
  NOR2X1 U546 ( .A(n802), .B(n1385), .Y(N182) );
  NOR4BX1 U547 ( .AN(n1381), .B(n707), .C(n1386), .D(n1387), .Y(n1385) );
  AOI2BB1X1 U548 ( .A0N(n1388), .A1N(n1389), .B0(n802), .Y(N181) );
  OAI2BB1X1 U549 ( .A0N(n1382), .A1N(n707), .B0(n1381), .Y(n1389) );
  MXI2X1 U550 ( .A(n13901), .B(n1391), .S0(n1392), .Y(n1381) );
  CLKINVX1 U551 ( .A(n1384), .Y(n1391) );
  NOR3X1 U552 ( .A(re_cs[0]), .B(re_cs[2]), .C(n942), .Y(n707) );
  OAI2BB2XL U553 ( .B0(n941), .B1(n1393), .A0N(n1387), .A1N(re_cs[0]), .Y(
        n1388) );
  OAI21XL U554 ( .A0(n1382), .A1(n1394), .B0(n1384), .Y(n1387) );
  NAND3X1 U555 ( .A(re_cs[2]), .B(n1395), .C(n941), .Y(n1384) );
  CLKINVX1 U556 ( .A(n1383), .Y(n1394) );
  XOR2X1 U557 ( .A(n1396), .B(re_cs[0]), .Y(n1393) );
  NAND2BX1 U558 ( .AN(N143), .B(n1187), .Y(N168) );
  NAND2BX1 U559 ( .AN(N141), .B(n1188), .Y(N166) );
  NAND2BX1 U560 ( .AN(N140), .B(n1187), .Y(N165) );
  NAND2BX1 U561 ( .AN(N139), .B(n1188), .Y(N164) );
  NAND2BX1 U562 ( .AN(N148), .B(n796), .Y(N163) );
  NAND2BX1 U563 ( .AN(N147), .B(n796), .Y(N162) );
  NAND2BX1 U564 ( .AN(N146), .B(n796), .Y(N161) );
  NAND2BX1 U565 ( .AN(N145), .B(n1187), .Y(N160) );
  AOI221XL U566 ( .A0(n1382), .A1(n1383), .B0(n1392), .B1(n13901), .C0(n1386), 
        .Y(n1397) );
  NOR3X1 U567 ( .A(n1396), .B(n941), .C(n1395), .Y(n1386) );
  MXI2X1 U568 ( .A(n1398), .B(n1399), .S0(re_cs[2]), .Y(n1396) );
  NOR2X1 U569 ( .A(n14001), .B(n1401), .Y(n1399) );
  NOR2X1 U570 ( .A(n1402), .B(n1403), .Y(n1398) );
  NOR2X1 U571 ( .A(n1401), .B(n1403), .Y(n1392) );
  NOR2X1 U572 ( .A(n14001), .B(n1402), .Y(n1382) );
  XOR2X1 U573 ( .A(n942), .B(write_addr_low[4]), .Y(n1258) );
  XOR2X1 U574 ( .A(n1243), .B(n941), .Y(n1261) );
  CLE_DW01_inc_0 add_249_S2 ( .A(index_cnt), .SUM({N343, N342, N341, N340, 
        N339, N338, N337, N336}) );
  CLE_DW01_inc_1 add_94 ( .A({write_addr_high, write_addr_low, N149, rw}), 
        .SUM({N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138}) );
  CLE_DW01_inc_2 add_83 ( .A({rom_a_high, rom_a_low, cnt[3:1], n1177}), .SUM({
        N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114}) );
  CLE_DW01_inc_3 add_76_S2 ( .A(times), .SUM({N88, N87, N86, N85, N84, N83, 
        N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, 
        N68}) );
  DFFQXL write_addr_high_reg_4_ ( .D(N163), .CK(clk), .Q(write_addr_high[4])
         );
  DFFQXL write_addr_low_reg_0_ ( .D(N164), .CK(clk), .Q(N149) );
  DFFX1 index_buffer_reg_28__7_ ( .D(n747), .CK(clk), .Q(index_buffer_28__7_), 
        .QN(n597) );
  DFFX1 index_buffer_reg_28__4_ ( .D(n7501), .CK(clk), .Q(index_buffer_28__4_), 
        .QN(n600) );
  DFFX1 index_buffer_reg_28__2_ ( .D(n752), .CK(clk), .Q(index_buffer_28__2_), 
        .QN(n602) );
  DFFX1 index_buffer_reg_28__1_ ( .D(n753), .CK(clk), .Q(index_buffer_28__1_), 
        .QN(n603) );
  DFFX1 index_buffer_reg_28__0_ ( .D(n754), .CK(clk), .Q(index_buffer_28__0_), 
        .QN(n604) );
  DFFX1 index_buffer_reg_29__6_ ( .D(n756), .CK(clk), .Q(index_buffer_29__6_), 
        .QN(n606) );
  DFFX1 index_buffer_reg_29__4_ ( .D(n758), .CK(clk), .Q(index_buffer_29__4_), 
        .QN(n608) );
  DFFX1 index_buffer_reg_29__2_ ( .D(n7601), .CK(clk), .Q(index_buffer_29__2_), 
        .QN(n610) );
  DFFX1 index_buffer_reg_29__0_ ( .D(n762), .CK(clk), .Q(index_buffer_29__0_), 
        .QN(n612) );
  EDFFTRX1 rd_buffer_reg_34_ ( .RN(n1437), .D(n242), .E(n1221), .CK(clk), .Q(
        n241) );
  EDFFTRX1 rd_buffer_reg_33_ ( .RN(n1438), .D(n243), .E(n1221), .CK(clk), .Q(
        n242) );
  EDFFTRX1 rd_buffer_reg_32_ ( .RN(n1437), .D(n244), .E(n1221), .CK(clk), .Q(
        n243) );
  EDFFTRX1 rd_buffer_reg_31_ ( .RN(n1438), .D(n245), .E(n1221), .CK(clk), .Q(
        n244) );
  EDFFTRX1 rd_buffer_reg_30_ ( .RN(n1437), .D(n246), .E(n1221), .CK(clk), .Q(
        n245) );
  EDFFTRX1 rd_buffer_reg_29_ ( .RN(n1438), .D(n247), .E(n1221), .CK(clk), .Q(
        n246) );
  EDFFTRX1 rd_buffer_reg_28_ ( .RN(n1437), .D(n248), .E(n1221), .CK(clk), .Q(
        n247) );
  EDFFTRX1 rd_buffer_reg_27_ ( .RN(n1438), .D(n249), .E(n1221), .CK(clk), .Q(
        n248) );
  EDFFTRX1 rd_buffer_reg_26_ ( .RN(n1437), .D(n250), .E(n1221), .CK(clk), .Q(
        n249) );
  EDFFTRX1 rd_buffer_reg_25_ ( .RN(n1438), .D(n251), .E(n1221), .CK(clk), .Q(
        n250) );
  EDFFTRX1 rd_buffer_reg_24_ ( .RN(n1437), .D(n252), .E(n1221), .CK(clk), .Q(
        n251) );
  EDFFTRX1 rd_buffer_reg_23_ ( .RN(n1438), .D(n253), .E(n1221), .CK(clk), .Q(
        n252) );
  EDFFTRX1 rd_buffer_reg_22_ ( .RN(n1437), .D(n254), .E(n1221), .CK(clk), .Q(
        n253) );
  EDFFTRX1 index_buffer_reg_27__0_ ( .RN(n1438), .D(index_buffer_28__0_), .E(
        n1221), .CK(clk), .Q(n234) );
  EDFFTRX1 index_buffer_reg_27__2_ ( .RN(n1437), .D(index_buffer_28__2_), .E(
        n1181), .CK(clk), .Q(n180) );
  EDFFTRX1 index_buffer_reg_27__1_ ( .RN(n1438), .D(index_buffer_28__1_), .E(
        n1183), .CK(clk), .Q(n207) );
  EDFFTRX1 index_buffer_reg_26__2_ ( .RN(n1437), .D(n180), .E(n1182), .CK(clk), 
        .Q(n179) );
  EDFFTRX1 index_buffer_reg_26__1_ ( .RN(n1438), .D(n207), .E(n1181), .CK(clk), 
        .Q(n206) );
  EDFFTRX1 index_buffer_reg_25__2_ ( .RN(n1437), .D(n179), .E(n1183), .CK(clk), 
        .Q(n178) );
  EDFFTRX1 index_buffer_reg_25__1_ ( .RN(n1438), .D(n206), .E(n1182), .CK(clk), 
        .Q(n205) );
  EDFFTRX1 index_buffer_reg_24__2_ ( .RN(n1437), .D(n178), .E(n1181), .CK(clk), 
        .Q(n177) );
  EDFFTRX1 index_buffer_reg_24__1_ ( .RN(n1437), .D(n205), .E(n1183), .CK(clk), 
        .Q(n204) );
  EDFFTRX1 index_buffer_reg_23__2_ ( .RN(n1438), .D(n177), .E(n1182), .CK(clk), 
        .Q(n176) );
  EDFFTRX1 index_buffer_reg_23__1_ ( .RN(n1437), .D(n204), .E(n1181), .CK(clk), 
        .Q(n203) );
  EDFFTRX1 index_buffer_reg_22__2_ ( .RN(n1437), .D(n176), .E(n1183), .CK(clk), 
        .Q(n175) );
  EDFFTRX1 index_buffer_reg_22__1_ ( .RN(n1438), .D(n203), .E(n1182), .CK(clk), 
        .Q(n202) );
  EDFFTRX1 index_buffer_reg_21__2_ ( .RN(n1437), .D(n175), .E(n1181), .CK(clk), 
        .Q(n174) );
  EDFFTRX1 index_buffer_reg_21__1_ ( .RN(n1437), .D(n202), .E(n1183), .CK(clk), 
        .Q(n201) );
  EDFFTRX1 index_buffer_reg_20__2_ ( .RN(n1438), .D(n174), .E(n1182), .CK(clk), 
        .Q(n173) );
  EDFFTRX1 index_buffer_reg_20__1_ ( .RN(n1437), .D(n201), .E(n1181), .CK(clk), 
        .Q(n200) );
  EDFFTRX1 index_buffer_reg_19__2_ ( .RN(n1437), .D(n173), .E(n1183), .CK(clk), 
        .Q(n172) );
  EDFFTRX1 index_buffer_reg_19__1_ ( .RN(n1438), .D(n200), .E(n1182), .CK(clk), 
        .Q(n199) );
  EDFFTRX1 index_buffer_reg_18__2_ ( .RN(n1437), .D(n172), .E(n1181), .CK(clk), 
        .Q(n171) );
  EDFFTRX1 index_buffer_reg_18__1_ ( .RN(n1437), .D(n199), .E(n1183), .CK(clk), 
        .Q(n198) );
  EDFFTRX1 index_buffer_reg_17__2_ ( .RN(n1438), .D(n171), .E(n1182), .CK(clk), 
        .Q(n170) );
  EDFFTRX1 index_buffer_reg_17__1_ ( .RN(n1437), .D(n198), .E(n1181), .CK(clk), 
        .Q(n197) );
  EDFFTRX1 index_buffer_reg_16__2_ ( .RN(n1437), .D(n170), .E(n1183), .CK(clk), 
        .Q(n169) );
  EDFFTRX1 index_buffer_reg_16__1_ ( .RN(n1438), .D(n197), .E(n1182), .CK(clk), 
        .Q(n196) );
  EDFFTRX1 index_buffer_reg_15__2_ ( .RN(n1437), .D(n169), .E(n1181), .CK(clk), 
        .Q(n1680) );
  EDFFTRX1 index_buffer_reg_15__1_ ( .RN(n1437), .D(n196), .E(n1183), .CK(clk), 
        .Q(n195) );
  EDFFTRX1 index_buffer_reg_14__2_ ( .RN(n1438), .D(n1680), .E(n1182), .CK(clk), .Q(n167) );
  EDFFTRX1 index_buffer_reg_14__1_ ( .RN(n1437), .D(n195), .E(n1181), .CK(clk), 
        .Q(n194) );
  EDFFTRX1 index_buffer_reg_13__1_ ( .RN(n1437), .D(n194), .E(n1182), .CK(clk), 
        .Q(n193) );
  EDFFTRX1 index_buffer_reg_13__0_ ( .RN(n1438), .D(n221), .E(n1181), .CK(clk), 
        .Q(n220) );
  EDFFTRX1 index_buffer_reg_12__1_ ( .RN(n1437), .D(n193), .E(n1183), .CK(clk), 
        .Q(n192) );
  EDFFTRX1 index_buffer_reg_12__0_ ( .RN(n1438), .D(n220), .E(n1182), .CK(clk), 
        .Q(n219) );
  EDFFTRX1 index_buffer_reg_11__1_ ( .RN(n1437), .D(n192), .E(n1181), .CK(clk), 
        .Q(n191) );
  EDFFTRX1 index_buffer_reg_11__0_ ( .RN(n1438), .D(n219), .E(n1183), .CK(clk), 
        .Q(n218) );
  EDFFTRX1 index_buffer_reg_10__1_ ( .RN(n1438), .D(n191), .E(n1182), .CK(clk), 
        .Q(n190) );
  EDFFTRX1 index_buffer_reg_10__0_ ( .RN(n1438), .D(n218), .E(n1181), .CK(clk), 
        .Q(n217) );
  EDFFTRX1 index_buffer_reg_9__1_ ( .RN(n1438), .D(n190), .E(n1183), .CK(clk), 
        .Q(n189) );
  EDFFTRX1 index_buffer_reg_9__0_ ( .RN(n1438), .D(n217), .E(n1182), .CK(clk), 
        .Q(n216) );
  EDFFTRX1 index_buffer_reg_8__1_ ( .RN(n1438), .D(n189), .E(n1181), .CK(clk), 
        .Q(n188) );
  EDFFTRX1 index_buffer_reg_8__0_ ( .RN(n1438), .D(n216), .E(n1183), .CK(clk), 
        .Q(n215) );
  EDFFTRX1 index_buffer_reg_7__1_ ( .RN(n1438), .D(n188), .E(n1182), .CK(clk), 
        .Q(n187) );
  EDFFTRX1 index_buffer_reg_7__0_ ( .RN(n1438), .D(n215), .E(n1181), .CK(clk), 
        .Q(n214) );
  EDFFTRX1 index_buffer_reg_6__1_ ( .RN(n1438), .D(n187), .E(n1183), .CK(clk), 
        .Q(n186) );
  EDFFTRX1 index_buffer_reg_6__0_ ( .RN(n1438), .D(n214), .E(n1182), .CK(clk), 
        .Q(n213) );
  EDFFTRX1 index_buffer_reg_5__1_ ( .RN(n1438), .D(n186), .E(n1181), .CK(clk), 
        .Q(n185) );
  EDFFTRX1 index_buffer_reg_5__0_ ( .RN(n1438), .D(n213), .E(n1183), .CK(clk), 
        .Q(n212) );
  EDFFTRX1 index_buffer_reg_4__1_ ( .RN(n1438), .D(n185), .E(n1182), .CK(clk), 
        .Q(n184) );
  EDFFTRX1 index_buffer_reg_4__0_ ( .RN(n1438), .D(n212), .E(n1181), .CK(clk), 
        .Q(n211) );
  EDFFTRX1 index_buffer_reg_3__1_ ( .RN(n1438), .D(n184), .E(n1183), .CK(clk), 
        .Q(n1830) );
  EDFFTRX1 index_buffer_reg_3__0_ ( .RN(n1438), .D(n211), .E(n1182), .CK(clk), 
        .Q(n210) );
  EDFFTRX1 index_buffer_reg_2__1_ ( .RN(n1438), .D(n1830), .E(n1181), .CK(clk), 
        .Q(n1820) );
  EDFFTRX1 index_buffer_reg_2__0_ ( .RN(n1438), .D(n210), .E(n1183), .CK(clk), 
        .Q(n209) );
  EDFFTRX1 index_buffer_reg_1__1_ ( .RN(n1438), .D(n1820), .E(n1182), .CK(clk), 
        .Q(n1810) );
  EDFFTRX1 index_buffer_reg_1__0_ ( .RN(n1438), .D(n209), .E(n1181), .CK(clk), 
        .Q(n208) );
  EDFFTRX1 rd_buffer_reg_21_ ( .RN(n1438), .D(n255), .E(n1221), .CK(clk), .Q(
        n254) );
  EDFFTRX1 rd_buffer_reg_20_ ( .RN(n1438), .D(n256), .E(n1221), .CK(clk), .Q(
        n255) );
  EDFFTRX1 rd_buffer_reg_19_ ( .RN(n1438), .D(n257), .E(n1221), .CK(clk), .Q(
        n256) );
  EDFFTRX1 rd_buffer_reg_18_ ( .RN(n1438), .D(n258), .E(n1221), .CK(clk), .Q(
        n257) );
  EDFFTRX1 rd_buffer_reg_17_ ( .RN(n1438), .D(n259), .E(n1221), .CK(clk), .Q(
        n258) );
  EDFFTRX1 rd_buffer_reg_16_ ( .RN(n1438), .D(n260), .E(n1221), .CK(clk), .Q(
        n259) );
  EDFFTRX1 rd_buffer_reg_15_ ( .RN(n1438), .D(n261), .E(n1221), .CK(clk), .Q(
        n260) );
  EDFFTRX1 rd_buffer_reg_14_ ( .RN(n1438), .D(n262), .E(n1221), .CK(clk), .Q(
        n261) );
  EDFFTRX1 rd_buffer_reg_13_ ( .RN(n1438), .D(rd_buffer[12]), .E(n1221), .CK(
        clk), .Q(n262) );
  EDFFTRX1 rd_buffer_reg_12_ ( .RN(n1438), .D(n263), .E(n1221), .CK(clk), .Q(
        rd_buffer[12]) );
  EDFFTRX1 rd_buffer_reg_11_ ( .RN(n1438), .D(n264), .E(n1221), .CK(clk), .Q(
        n263) );
  EDFFTRX1 rd_buffer_reg_10_ ( .RN(n1438), .D(n265), .E(n1221), .CK(clk), .Q(
        n264) );
  EDFFTRX1 rd_buffer_reg_9_ ( .RN(n1438), .D(rd_buffer[8]), .E(n1221), .CK(clk), .Q(n265) );
  EDFFTRX1 index_buffer_reg_26__0_ ( .RN(n1438), .D(n234), .E(n1221), .CK(clk), 
        .Q(n233) );
  EDFFTRX1 index_buffer_reg_25__0_ ( .RN(n1438), .D(n233), .E(n1221), .CK(clk), 
        .Q(n232) );
  EDFFTRX1 index_buffer_reg_24__0_ ( .RN(n1438), .D(n232), .E(n1221), .CK(clk), 
        .Q(n231) );
  EDFFTRX1 index_buffer_reg_23__0_ ( .RN(n1438), .D(n231), .E(n1221), .CK(clk), 
        .Q(n230) );
  EDFFTRX1 index_buffer_reg_22__0_ ( .RN(n1438), .D(n230), .E(n1221), .CK(clk), 
        .Q(n229) );
  EDFFTRX1 index_buffer_reg_21__0_ ( .RN(n1438), .D(n229), .E(n1221), .CK(clk), 
        .Q(n228) );
  EDFFTRX1 index_buffer_reg_20__0_ ( .RN(n1438), .D(n228), .E(n1221), .CK(clk), 
        .Q(n227) );
  EDFFTRX1 index_buffer_reg_19__0_ ( .RN(n1438), .D(n227), .E(n1221), .CK(clk), 
        .Q(n226) );
  EDFFTRX1 index_buffer_reg_18__0_ ( .RN(n1438), .D(n226), .E(n1221), .CK(clk), 
        .Q(n225) );
  EDFFTRX1 index_buffer_reg_17__0_ ( .RN(n1438), .D(n225), .E(n1221), .CK(clk), 
        .Q(n224) );
  EDFFTRX1 index_buffer_reg_16__0_ ( .RN(n1438), .D(n224), .E(n1221), .CK(clk), 
        .Q(n223) );
  EDFFTRX1 index_buffer_reg_15__0_ ( .RN(n1438), .D(n223), .E(n1221), .CK(clk), 
        .Q(n222) );
  EDFFTRX1 index_buffer_reg_14__0_ ( .RN(n1438), .D(n222), .E(n1221), .CK(clk), 
        .Q(n221) );
  EDFFTRX1 index_buffer_reg_7__3_ ( .RN(n1438), .D(n26), .E(n1183), .CK(clk), 
        .Q(n25) );
  EDFFTRX1 index_buffer_reg_6__3_ ( .RN(n1438), .D(n25), .E(n12201), .CK(clk), 
        .Q(n24) );
  EDFFTRX1 index_buffer_reg_5__3_ ( .RN(n1437), .D(n24), .E(n1177), .CK(clk), 
        .Q(n23) );
  EDFFTRX1 index_buffer_reg_4__3_ ( .RN(n1437), .D(n23), .E(n1181), .CK(clk), 
        .Q(n22) );
  EDFFTRX1 index_buffer_reg_4__2_ ( .RN(n1438), .D(n1580), .E(n1183), .CK(clk), 
        .Q(n1570) );
  EDFFTRX1 index_buffer_reg_3__3_ ( .RN(n1438), .D(n22), .E(n1219), .CK(clk), 
        .Q(n21) );
  EDFFTRX1 index_buffer_reg_2__3_ ( .RN(n1438), .D(n21), .E(n1177), .CK(clk), 
        .Q(n20) );
  EDFFTRX1 index_buffer_reg_27__5_ ( .RN(n14101), .D(index_buffer_28__5_), .E(
        n1178), .CK(clk), .Q(n99) );
  EDFFTRX1 index_buffer_reg_27__4_ ( .RN(n14101), .D(index_buffer_28__4_), .E(
        n1221), .CK(clk), .Q(n720) );
  EDFFTRX1 index_buffer_reg_27__3_ ( .RN(n14101), .D(index_buffer_28__3_), .E(
        n1182), .CK(clk), .Q(n45) );
  EDFFTRX1 index_buffer_reg_26__5_ ( .RN(n14101), .D(n99), .E(n1179), .CK(clk), 
        .Q(n98) );
  EDFFTRX1 index_buffer_reg_26__4_ ( .RN(n14101), .D(n720), .E(n12201), .CK(
        clk), .Q(n710) );
  EDFFTRX1 index_buffer_reg_26__3_ ( .RN(n14101), .D(n45), .E(n1177), .CK(clk), 
        .Q(n44) );
  EDFFTRX1 index_buffer_reg_25__5_ ( .RN(n14101), .D(n98), .E(n11801), .CK(clk), .Q(n97) );
  EDFFTRX1 index_buffer_reg_25__4_ ( .RN(n14101), .D(n710), .E(n1177), .CK(clk), .Q(n700) );
  EDFFTRX1 index_buffer_reg_25__3_ ( .RN(n14101), .D(n44), .E(n1221), .CK(clk), 
        .Q(n43) );
  EDFFTRX1 index_buffer_reg_24__5_ ( .RN(n14101), .D(n97), .E(n1178), .CK(clk), 
        .Q(n96) );
  EDFFTRX1 index_buffer_reg_24__4_ ( .RN(n14101), .D(n700), .E(n1221), .CK(clk), .Q(n690) );
  EDFFTRX1 index_buffer_reg_24__3_ ( .RN(n14101), .D(n43), .E(n12201), .CK(clk), .Q(n42) );
  EDFFTRX1 index_buffer_reg_23__5_ ( .RN(n14101), .D(n96), .E(n1179), .CK(clk), 
        .Q(n95) );
  EDFFTRX1 index_buffer_reg_23__4_ ( .RN(n14101), .D(n690), .E(n12201), .CK(
        clk), .Q(n680) );
  EDFFTRX1 index_buffer_reg_23__3_ ( .RN(n14101), .D(n42), .E(n1177), .CK(clk), 
        .Q(n41) );
  EDFFTRX1 index_buffer_reg_22__5_ ( .RN(n14101), .D(n95), .E(n11801), .CK(clk), .Q(n94) );
  EDFFTRX1 index_buffer_reg_22__4_ ( .RN(n14101), .D(n680), .E(n1177), .CK(clk), .Q(n67) );
  EDFFTRX1 index_buffer_reg_22__3_ ( .RN(n14101), .D(n41), .E(n1221), .CK(clk), 
        .Q(n40) );
  EDFFTRX1 index_buffer_reg_21__5_ ( .RN(n14101), .D(n94), .E(n1178), .CK(clk), 
        .Q(n93) );
  EDFFTRX1 index_buffer_reg_21__4_ ( .RN(n14101), .D(n67), .E(n1221), .CK(clk), 
        .Q(n66) );
  EDFFTRX1 index_buffer_reg_21__3_ ( .RN(n14101), .D(n40), .E(cnt[0]), .CK(clk), .Q(n39) );
  EDFFTRX1 index_buffer_reg_20__5_ ( .RN(n14101), .D(n93), .E(n1179), .CK(clk), 
        .Q(n92) );
  EDFFTRX1 index_buffer_reg_20__4_ ( .RN(n14101), .D(n66), .E(n12201), .CK(clk), .Q(n65) );
  EDFFTRX1 index_buffer_reg_20__3_ ( .RN(n14101), .D(n39), .E(n1177), .CK(clk), 
        .Q(n38) );
  EDFFTRX1 index_buffer_reg_19__5_ ( .RN(n14101), .D(n92), .E(n11801), .CK(clk), .Q(n91) );
  EDFFTRX1 index_buffer_reg_19__4_ ( .RN(n14101), .D(n65), .E(n1177), .CK(clk), 
        .Q(n64) );
  EDFFTRX1 index_buffer_reg_19__3_ ( .RN(n14101), .D(n38), .E(n1179), .CK(clk), 
        .Q(n37) );
  EDFFTRX2 index_buffer_reg_0__2_ ( .RN(n1196), .D(n1540), .E(cnt[0]), .CK(clk), .Q(n1567), .QN(n1308) );
  DFFX2 re_cs_reg_2_ ( .D(N183), .CK(clk), .Q(re_cs[2]), .QN(n1257) );
  DFFX2 re_cs_reg_1_ ( .D(N182), .CK(clk), .Q(n941), .QN(n942) );
  DFFX2 cs_reg ( .D(n787), .CK(clk), .Q(cs), .QN(n1412) );
  DFFQX1 rd_buffer_reg_7_ ( .D(n788), .CK(clk), .Q(rd_buffer[7]) );
  DFFQX1 write_addr_high_reg_3_ ( .D(N162), .CK(clk), .Q(write_addr_high[3])
         );
  DFFQX1 write_addr_high_reg_2_ ( .D(N161), .CK(clk), .Q(write_addr_high[2])
         );
  DFFQX1 write_addr_low_reg_2_ ( .D(N166), .CK(clk), .Q(write_addr_low[2]) );
  DFFQX1 write_addr_high_reg_1_ ( .D(N160), .CK(clk), .Q(write_addr_high[1])
         );
  DFFQX1 write_addr_low_reg_4_ ( .D(N168), .CK(clk), .Q(write_addr_low[4]) );
  NOR3X1 U234 ( .A(n942), .B(re_cs[2]), .C(n1395), .Y(n1383) );
  INVXL U260 ( .A(n1567), .Y(n14341) );
  INVX12 U264 ( .A(n14341), .Y(sram_d[2]) );
  CLKBUFX3 U345 ( .A(n14101), .Y(n1189) );
  INVX4 U347 ( .A(n802), .Y(n14101) );
  CLKINVX6 U349 ( .A(n1189), .Y(n1436) );
  INVX12 U351 ( .A(n1436), .Y(n1437) );
  INVX16 U537 ( .A(n1436), .Y(n1438) );
endmodule

